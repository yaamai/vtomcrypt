module tomcrypt

#include "@VMODROOT/tc_helper_top.h"

#flag -I @VMODROOT/tommath
#flag @VMODROOT/libtommath/bn_cutoffs.o
#flag @VMODROOT/libtommath/bn_deprecated.o
#flag @VMODROOT/libtommath/bn_mp_2expt.o
#flag @VMODROOT/libtommath/bn_mp_abs.o
#flag @VMODROOT/libtommath/bn_mp_add.o
#flag @VMODROOT/libtommath/bn_mp_add_d.o
#flag @VMODROOT/libtommath/bn_mp_addmod.o
#flag @VMODROOT/libtommath/bn_mp_and.o
#flag @VMODROOT/libtommath/bn_mp_clamp.o
#flag @VMODROOT/libtommath/bn_mp_clear.o
#flag @VMODROOT/libtommath/bn_mp_clear_multi.o
#flag @VMODROOT/libtommath/bn_mp_cmp.o
#flag @VMODROOT/libtommath/bn_mp_cmp_d.o
#flag @VMODROOT/libtommath/bn_mp_cmp_mag.o
#flag @VMODROOT/libtommath/bn_mp_cnt_lsb.o
#flag @VMODROOT/libtommath/bn_mp_complement.o
#flag @VMODROOT/libtommath/bn_mp_copy.o
#flag @VMODROOT/libtommath/bn_mp_count_bits.o
#flag @VMODROOT/libtommath/bn_mp_decr.o
#flag @VMODROOT/libtommath/bn_mp_div.o
#flag @VMODROOT/libtommath/bn_mp_div_2.o
#flag @VMODROOT/libtommath/bn_mp_div_2d.o
#flag @VMODROOT/libtommath/bn_mp_div_3.o
#flag @VMODROOT/libtommath/bn_mp_div_d.o
#flag @VMODROOT/libtommath/bn_mp_dr_is_modulus.o
#flag @VMODROOT/libtommath/bn_mp_dr_reduce.o
#flag @VMODROOT/libtommath/bn_mp_dr_setup.o
#flag @VMODROOT/libtommath/bn_mp_error_to_string.o
#flag @VMODROOT/libtommath/bn_mp_exch.o
#flag @VMODROOT/libtommath/bn_mp_expt_u32.o
#flag @VMODROOT/libtommath/bn_mp_exptmod.o
#flag @VMODROOT/libtommath/bn_mp_exteuclid.o
#flag @VMODROOT/libtommath/bn_mp_fread.o
#flag @VMODROOT/libtommath/bn_mp_from_sbin.o
#flag @VMODROOT/libtommath/bn_mp_from_ubin.o
#flag @VMODROOT/libtommath/bn_mp_fwrite.o
#flag @VMODROOT/libtommath/bn_mp_gcd.o
#flag @VMODROOT/libtommath/bn_mp_get_double.o
#flag @VMODROOT/libtommath/bn_mp_get_i32.o
#flag @VMODROOT/libtommath/bn_mp_get_i64.o
#flag @VMODROOT/libtommath/bn_mp_get_l.o
#flag @VMODROOT/libtommath/bn_mp_get_ll.o
#flag @VMODROOT/libtommath/bn_mp_get_mag_u32.o
#flag @VMODROOT/libtommath/bn_mp_get_mag_u64.o
#flag @VMODROOT/libtommath/bn_mp_get_mag_ul.o
#flag @VMODROOT/libtommath/bn_mp_get_mag_ull.o
#flag @VMODROOT/libtommath/bn_mp_grow.o
#flag @VMODROOT/libtommath/bn_mp_incr.o
#flag @VMODROOT/libtommath/bn_mp_init.o
#flag @VMODROOT/libtommath/bn_mp_init_copy.o
#flag @VMODROOT/libtommath/bn_mp_init_i32.o
#flag @VMODROOT/libtommath/bn_mp_init_i64.o
#flag @VMODROOT/libtommath/bn_mp_init_l.o
#flag @VMODROOT/libtommath/bn_mp_init_ll.o
#flag @VMODROOT/libtommath/bn_mp_init_multi.o
#flag @VMODROOT/libtommath/bn_mp_init_set.o
#flag @VMODROOT/libtommath/bn_mp_init_size.o
#flag @VMODROOT/libtommath/bn_mp_init_u32.o
#flag @VMODROOT/libtommath/bn_mp_init_u64.o
#flag @VMODROOT/libtommath/bn_mp_init_ul.o
#flag @VMODROOT/libtommath/bn_mp_init_ull.o
#flag @VMODROOT/libtommath/bn_mp_invmod.o
#flag @VMODROOT/libtommath/bn_mp_is_square.o
#flag @VMODROOT/libtommath/bn_mp_iseven.o
#flag @VMODROOT/libtommath/bn_mp_isodd.o
#flag @VMODROOT/libtommath/bn_mp_kronecker.o
#flag @VMODROOT/libtommath/bn_mp_lcm.o
#flag @VMODROOT/libtommath/bn_mp_log_u32.o
#flag @VMODROOT/libtommath/bn_mp_lshd.o
#flag @VMODROOT/libtommath/bn_mp_mod.o
#flag @VMODROOT/libtommath/bn_mp_mod_2d.o
#flag @VMODROOT/libtommath/bn_mp_mod_d.o
#flag @VMODROOT/libtommath/bn_mp_montgomery_calc_normalization.o
#flag @VMODROOT/libtommath/bn_mp_montgomery_reduce.o
#flag @VMODROOT/libtommath/bn_mp_montgomery_setup.o
#flag @VMODROOT/libtommath/bn_mp_mul.o
#flag @VMODROOT/libtommath/bn_mp_mul_2.o
#flag @VMODROOT/libtommath/bn_mp_mul_2d.o
#flag @VMODROOT/libtommath/bn_mp_mul_d.o
#flag @VMODROOT/libtommath/bn_mp_mulmod.o
#flag @VMODROOT/libtommath/bn_mp_neg.o
#flag @VMODROOT/libtommath/bn_mp_or.o
#flag @VMODROOT/libtommath/bn_mp_pack.o
#flag @VMODROOT/libtommath/bn_mp_pack_count.o
#flag @VMODROOT/libtommath/bn_mp_prime_fermat.o
#flag @VMODROOT/libtommath/bn_mp_prime_frobenius_underwood.o
#flag @VMODROOT/libtommath/bn_mp_prime_is_prime.o
#flag @VMODROOT/libtommath/bn_mp_prime_miller_rabin.o
#flag @VMODROOT/libtommath/bn_mp_prime_next_prime.o
#flag @VMODROOT/libtommath/bn_mp_prime_rabin_miller_trials.o
#flag @VMODROOT/libtommath/bn_mp_prime_rand.o
#flag @VMODROOT/libtommath/bn_mp_prime_strong_lucas_selfridge.o
#flag @VMODROOT/libtommath/bn_mp_radix_size.o
#flag @VMODROOT/libtommath/bn_mp_radix_smap.o
#flag @VMODROOT/libtommath/bn_mp_rand.o
#flag @VMODROOT/libtommath/bn_mp_read_radix.o
#flag @VMODROOT/libtommath/bn_mp_reduce.o
#flag @VMODROOT/libtommath/bn_mp_reduce_2k.o
#flag @VMODROOT/libtommath/bn_mp_reduce_2k_l.o
#flag @VMODROOT/libtommath/bn_mp_reduce_2k_setup.o
#flag @VMODROOT/libtommath/bn_mp_reduce_2k_setup_l.o
#flag @VMODROOT/libtommath/bn_mp_reduce_is_2k.o
#flag @VMODROOT/libtommath/bn_mp_reduce_is_2k_l.o
#flag @VMODROOT/libtommath/bn_mp_reduce_setup.o
#flag @VMODROOT/libtommath/bn_mp_root_u32.o
#flag @VMODROOT/libtommath/bn_mp_rshd.o
#flag @VMODROOT/libtommath/bn_mp_sbin_size.o
#flag @VMODROOT/libtommath/bn_mp_set.o
#flag @VMODROOT/libtommath/bn_mp_set_double.o
#flag @VMODROOT/libtommath/bn_mp_set_i32.o
#flag @VMODROOT/libtommath/bn_mp_set_i64.o
#flag @VMODROOT/libtommath/bn_mp_set_l.o
#flag @VMODROOT/libtommath/bn_mp_set_ll.o
#flag @VMODROOT/libtommath/bn_mp_set_u32.o
#flag @VMODROOT/libtommath/bn_mp_set_u64.o
#flag @VMODROOT/libtommath/bn_mp_set_ul.o
#flag @VMODROOT/libtommath/bn_mp_set_ull.o
#flag @VMODROOT/libtommath/bn_mp_shrink.o
#flag @VMODROOT/libtommath/bn_mp_signed_rsh.o
#flag @VMODROOT/libtommath/bn_mp_sqr.o
#flag @VMODROOT/libtommath/bn_mp_sqrmod.o
#flag @VMODROOT/libtommath/bn_mp_sqrt.o
#flag @VMODROOT/libtommath/bn_mp_sqrtmod_prime.o
#flag @VMODROOT/libtommath/bn_mp_sub.o
#flag @VMODROOT/libtommath/bn_mp_sub_d.o
#flag @VMODROOT/libtommath/bn_mp_submod.o
#flag @VMODROOT/libtommath/bn_mp_to_radix.o
#flag @VMODROOT/libtommath/bn_mp_to_sbin.o
#flag @VMODROOT/libtommath/bn_mp_to_ubin.o
#flag @VMODROOT/libtommath/bn_mp_ubin_size.o
#flag @VMODROOT/libtommath/bn_mp_unpack.o
#flag @VMODROOT/libtommath/bn_mp_xor.o
#flag @VMODROOT/libtommath/bn_mp_zero.o
#flag @VMODROOT/libtommath/bn_prime_tab.o
#flag @VMODROOT/libtommath/bn_s_mp_add.o
#flag @VMODROOT/libtommath/bn_s_mp_balance_mul.o
#flag @VMODROOT/libtommath/bn_s_mp_exptmod.o
#flag @VMODROOT/libtommath/bn_s_mp_exptmod_fast.o
#flag @VMODROOT/libtommath/bn_s_mp_get_bit.o
#flag @VMODROOT/libtommath/bn_s_mp_invmod_fast.o
#flag @VMODROOT/libtommath/bn_s_mp_invmod_slow.o
#flag @VMODROOT/libtommath/bn_s_mp_karatsuba_mul.o
#flag @VMODROOT/libtommath/bn_s_mp_karatsuba_sqr.o
#flag @VMODROOT/libtommath/bn_s_mp_montgomery_reduce_fast.o
#flag @VMODROOT/libtommath/bn_s_mp_mul_digs.o
#flag @VMODROOT/libtommath/bn_s_mp_mul_digs_fast.o
#flag @VMODROOT/libtommath/bn_s_mp_mul_high_digs.o
#flag @VMODROOT/libtommath/bn_s_mp_mul_high_digs_fast.o
#flag @VMODROOT/libtommath/bn_s_mp_prime_is_divisible.o
#flag @VMODROOT/libtommath/bn_s_mp_rand_jenkins.o
#flag @VMODROOT/libtommath/bn_s_mp_rand_platform.o
#flag @VMODROOT/libtommath/bn_s_mp_reverse.o
#flag @VMODROOT/libtommath/bn_s_mp_sqr.o
#flag @VMODROOT/libtommath/bn_s_mp_sqr_fast.o
#flag @VMODROOT/libtommath/bn_s_mp_sub.o
#flag @VMODROOT/libtommath/bn_s_mp_toom_mul.o
#flag @VMODROOT/libtommath/bn_s_mp_toom_sqr.o